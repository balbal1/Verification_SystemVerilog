module FSM_tb(FSM_if.TEST _if);
    
    initial begin
    
        $stop;
    end
    
endmodule

module FSM_monitor (FSM_if.MONITOR _if);
    
    initial begin
        $monitor("");
    end
    
endmodule

module FSM(FSM_if.DUT _if);
    
endmodule

module counter_monitor (counter_if.MONITOR _if);
    
    initial begin
        $monitor("");
    end
    
endmodule

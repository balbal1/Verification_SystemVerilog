module FSM_sva (FSM_if.DUT _if);
    
endmodule
